module core

import quickjs
