module core

pub fn test() {
	println('Hello from V')
}
